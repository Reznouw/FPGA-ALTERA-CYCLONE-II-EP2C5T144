library verilog;
use verilog.vl_types.all;
entity ejem_vlg_vec_tst is
end ejem_vlg_vec_tst;
