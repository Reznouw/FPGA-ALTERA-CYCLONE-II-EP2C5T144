library verilog;
use verilog.vl_types.all;
entity TF2_vlg_vec_tst is
end TF2_vlg_vec_tst;
