library verilog;
use verilog.vl_types.all;
entity labcalificado1_vlg_vec_tst is
end labcalificado1_vlg_vec_tst;
