library verilog;
use verilog.vl_types.all;
entity labcalificado1_vlg_check_tst is
    port(
        data_out        : in     vl_logic_vector(4 downto 0);
        sampler_rx      : in     vl_logic
    );
end labcalificado1_vlg_check_tst;
